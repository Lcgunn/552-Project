			//this determines if the alu gets imm or reg
module control_logic(input [3:0]Instr, output imm_or_reg);
	

endmodule
