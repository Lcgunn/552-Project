module cpu (output hlt, output pc[15:0], input clk, input rst_n);
	
endmodule